`timescale 1ns / 1ps

//========================================================================================================================
//                                                     Description
//========================================================================================================================
/*

Engineer   : HammerMeow
Date       : 07.07.2025 | 23:17

Description: lorem ipsum

*/
//========================================================================================================================

module test_module_tb;

//========================================================================================================================
//                                                  Parameters of UUT
//========================================================================================================================

parameter DATA_W = 8;

//========================================================================================================================
//                                                        Inputs
//========================================================================================================================

reg                     clk_in;
reg                     reset_in;

reg [(DATA_W-1):0]      data_in;

wire [(DATA_W-1):0]     out_0;
wire                    out_valid_0;
wire [(DATA_W-1):0]     out_1;
wire                    out_valid_1;
wire [(DATA_W-1):0]     out_2;
wire                    out_valid_2;
wire [(DATA_W-1):0]     out_3;
wire                    out_valid_3;

//========================================================================================================================
//                                                       Outputs
//========================================================================================================================



//========================================================================================================================
//                                              Parameters for simulation
//========================================================================================================================

parameter PERIOD = 10;
parameter DATA_FROM_EXAMPLE = 4;

//========================================================================================================================
//                                               Vars and genvar signals
//========================================================================================================================

integer en_display = 0;
integer cnt = 0;

//========================================================================================================================
//                                                       Includes
//========================================================================================================================



//========================================================================================================================
//                                                         UUT
//========================================================================================================================

test_module
#(
    .DATA_W(DATA_W)
) uut (
    .clk_in(clk_in),
    .reset_in(reset_in),
    .data_in(data_in),
    .out_0(out_0),
    .out_valid_0(out_valid_0),
    .out_1(out_1),
    .out_valid_1(out_valid_1),
    .out_2(out_2),
    .out_valid_2(out_valid_2),
    .out_3(out_3),
    .out_valid_3(out_valid_3)
);

//========================================================================================================================
//                                                       Initial
//========================================================================================================================

initial begin
    data_in  = 0;
    reset_in = 1;
    #(PERIOD/2);
    #(PERIOD*15);
    reset_in = 0;
    #(PERIOD*20);
    #(PERIOD/2);

    // user code
    if (DATA_FROM_EXAMPLE == 1) begin
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd2;
        #(PERIOD);
        en_display = 1;
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd2;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd2;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD*2);
        en_display = 0;
    end

    if (DATA_FROM_EXAMPLE == 2) begin
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd2;
        #(PERIOD);
        en_display = 1;
        data_in <= 8'd3;
        #(PERIOD);
        data_in <= 8'd4;
        #(PERIOD);
        data_in <= 8'd3;
        #(PERIOD);
        data_in <= 8'd2;
        #(PERIOD);
        data_in <= 8'd3;
        #(PERIOD);
        data_in <= 8'd4;
        #(PERIOD);
        data_in <= 8'd3;
        #(PERIOD);
        data_in <= 8'd4;
        #(PERIOD*2);
        en_display = 0;
    end

    if (DATA_FROM_EXAMPLE == 3) begin
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD);
        en_display = 1;
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD);
        data_in <= 8'd1;
        #(PERIOD*2);
        en_display = 0;
    end

    if (DATA_FROM_EXAMPLE == 4) begin
        data_in <= 8'd0;
        #(PERIOD);
        data_in <= 8'd0;
        #(PERIOD);
        en_display = 1;
        data_in <= 8'd0;
        #(PERIOD);
        data_in <= 8'd0;
        #(PERIOD);
        data_in <= 8'd0;
        #(PERIOD);
        data_in <= 8'd0;
        #(PERIOD);
        data_in <= 8'd0;
        #(PERIOD*2);
        en_display = 0;
    end
end

//========================================================================================================================
//                                                    Support logic
//========================================================================================================================

always @(posedge clk_in) begin
    if (en_display == 1) begin
        $display("num %d: out_0 = %h | out_1 = %h | out_2 = %h | out_3 = %h;", cnt, out_0, out_1, out_2, out_3);
        cnt = cnt + 1;
    end
end

always begin
    clk_in = 1'b1;
    #(PERIOD/2);
    clk_in = 1'b0;
    #(PERIOD/2);
end

//========================================================================================================================
//                                                     Local tasks
//========================================================================================================================



endmodule
